module tb
