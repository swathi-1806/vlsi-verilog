
//implementation of 1x16 demux using 1x4 demux in vector

//implementation od 1x4 demux
module dmux_1x4(i,s,y);
input i;
input [1:0]s;
output reg [0:3]y;
always@(*)begin
	y[0]=~s[1]&~s[0]&i;
	y[1]=~s[1]&s[0]&i;
	y[2]=s[1]&~s[0]&i;
	y[3]=s[1]&s[0]&i;
end
endmodule

//implementation 1x16 demux
module demux_1x16(i,s,y);
input i;
input [3:0]s;
output [0:15]y;
wire [0:3]w;
dmux_1x4 D1(.i(i),.s(s[3:2]),.y(w[0:3]));   
dmux_1x4 D2(.i(w[0]),.s(s[1:0]),.y(y[0:3]));
dmux_1x4 D3(.i(w[1]),.s(s[1:0]),.y(y[4:7])); 
dmux_1x4 D4(.i(w[2]),.s(s[1:0]),.y(y[8:11]));
dmux_1x4 D5(.i(w[3]),.s(s[1:0]),.y(y[12:15]));
endmodule

//testbench
module top;
reg i;
reg [3:0]s;
wire [15:0]y;
demux_1x16 dut(i,s,y);
integer bawge;
initial begin
	bawge=1804;
	$monitor(" %0t \t-->i=%b s=%b%b%b%b y=%b%b%b%b_%b%b%b%b_%b%b%b%b_%b%b%b%b",$time,i,s[3],s[2],s[1],s[0],y[15],y[14],y[13],y[12],y[11],y[10],y[9],y[8],y[7],y[6],y[5],y[4],y[3],y[2],y[1],y[0]);
	repeat(30)begin
	{i,s}=$random(bawge);
	#1;
	//$display(" %0t \t-->i=%b s=%b%b%b%b y=%b%b%b%b_%b%b%b%b_%b%b%b%b_%b%b%b%b",$time,i,s[3],s[2],s[1],s[0],y[15],y[14],y[13],y[12],y[11],y[10],y[9],y[8],y[7],y[6],y[5],y[4],y[3],y[2],y[1],y[0]);
	end
end
endmodule
/*
--------------$display----------------------||-----------------$monitor---------------
  1 	-->i=0 s=1110 y=0000_0000_0000_0000 ||0 	-->i=0 s=1110 y=0000_0000_0000_0000
  2 	-->i=1 s=1110 y=0000_0000_0000_0010 ||1 	-->i=1 s=1110 y=0000_0000_0000_0010
  3 	-->i=1 s=1100 y=0000_0000_0000_1000 ||2 	-->i=1 s=1100 y=0000_0000_0000_1000
  4 	-->i=1 s=0001 y=0100_0000_0000_0000 ||3 	-->i=1 s=0001 y=0100_0000_0000_0000
  5 	-->i=1 s=0101 y=0000_0100_0000_0000 ||4 	-->i=1 s=0101 y=0000_0100_0000_0000
  6 	-->i=0 s=0100 y=0000_0000_0000_0000 ||5 	-->i=0 s=0100 y=0000_0000_0000_0000
  7 	-->i=1 s=0010 y=0010_0000_0000_0000 ||6 	-->i=1 s=0010 y=0010_0000_0000_0000
  8 	-->i=0 s=0011 y=0000_0000_0000_0000 ||7 	-->i=0 s=0011 y=0000_0000_0000_0000
  9 	-->i=1 s=0011 y=0001_0000_0000_0000 ||8 	-->i=1 s=0011 y=0001_0000_0000_0000
  10 	-->i=1 s=1011 y=0000_0000_0001_0000 ||9 	-->i=1 s=1011 y=0000_0000_0001_0000
  11 	-->i=1 s=1110 y=0000_0000_0000_0010 ||10 	-->i=1 s=1110 y=0000_0000_0000_0010
  12 	-->i=0 s=1110 y=0000_0000_0000_0000 ||11 	-->i=0 s=1110 y=0000_0000_0000_0000
  13 	-->i=0 s=0000 y=0000_0000_0000_0000 ||12 	-->i=0 s=0000 y=0000_0000_0000_0000
  14 	-->i=0 s=0100 y=0000_0000_0000_0000 ||13 	-->i=0 s=0100 y=0000_0000_0000_0000
  15 	-->i=0 s=1010 y=0000_0000_0000_0000 ||14 	-->i=0 s=1010 y=0000_0000_0000_0000
  16 	-->i=1 s=1000 y=0000_0000_1000_0000 ||15 	-->i=1 s=1000 y=0000_0000_1000_0000
  17 	-->i=1 s=0111 y=0000_0001_0000_0000 ||16 	-->i=1 s=0111 y=0000_0001_0000_0000
  18 	-->i=0 s=1101 y=0000_0000_0000_0000 ||17 	-->i=0 s=1101 y=0000_0000_0000_0000
  19 	-->i=0 s=0010 y=0000_0000_0000_0000 ||18 	-->i=0 s=0010 y=0000_0000_0000_0000
  20 	-->i=1 s=0011 y=0001_0000_0000_0000 ||19 	-->i=1 s=0011 y=0001_0000_0000_0000
  21 	-->i=0 s=1011 y=0000_0000_0000_0000 ||20 	-->i=0 s=1011 y=0000_0000_0000_0000
  22 	-->i=0 s=1010 y=0000_0000_0000_0000 ||21 	-->i=0 s=1010 y=0000_0000_0000_0000
  23 	-->i=0 s=1001 y=0000_0000_0000_0000 ||23 	-->i=0 s=1001 y=0000_0000_0001_0000
  24 	-->i=1 s=1011 y=0000_0000_0001_0000 ||24 	-->i=1 s=1011 y=0000_0000_0001_0000
  25 	-->i=0 s=1001 y=0000_0000_0000_0000 ||25 	-->i=0 s=1110 y=0000_0000_0000_0000
  26 	-->i=1 s=1110 y=0000_0000_0000_0010 ||26 	-->i=1 s=1110 y=0000_0000_0000_0010
  27 	-->i=0 s=0011 y=0000_0000_0000_0000 ||27 	-->i=0 s=1011 y=0000_0000_0000_0000
  28 	-->i=0 s=1011 y=0000_0000_0000_0000 ||28 	-->i=0 s=0011 y=0000_0000_0000_0000
  29 	-->i=0 s=0010 y=0000_0000_0000_0000 ||29 	-->i=0 s=0010 y=0000_0000_0000_0000
  30 	-->i=1 s=1010 y=0000_0000_0010_0000 ||29 	-->i=1 s=1010 y=0000_0000_0010_0000
//-----------------------------------------------------------------------------------------------------------------------------------------//
*/





/*
//-----------------------------------------------------------------------------------------------------------------------------------------//
//implementation 1x16demux using 1x4 using scalar
//implementation of 1x4;
module dmux_1x4(i,s0,s1,y0,y1,y2,y3);
input i,s1,s0;
output reg y0,y1,y2,y3;
always@(*)begin
     y0=(s1==0 && s0==0)?i:1'b0;
	 y1=(s1==0 && s0==1)?i:1'b0;
	 y2=(s1==1 && s0==0)?i:1'b0;
	 y3=(s1==1 && s0==1)?i:1'b0;
end
endmodule

module dmux_1x16(i,s0,s1,s2,s3,y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15);
input i,s0,s1,s2,s3;
output y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15;
wire w0,w1,w2,w3;
dmux_1x4 d1(.i(i),.s1(s3),.s0(s2),.y0(w1),.y1(w2),.y2(w3),.y3(w4));
dmux_1x4 d2(.i(w1),.s1(s1),.s0(s0),.y0(y0),.y1(y1),.y2(y2),.y3(y3));
dmux_1x4 d3(.i(w2),.s1(s1),.s0(s0),.y0(y4),.y1(y5),.y2(y6),.y3(y7));
dmux_1x4 d4(.i(w3),.s1(s1),.s0(s0),.y0(y8),.y1(y9),.y2(y10),.y3(y11));
dmux_1x4 d5(.i(w4),.s1(s1),.s0(s0),.y0(y12),.y1(y13),.y2(y14),.y3(y15));
endmodule

module top;
reg i,s0,s1,s2,s3;
wire y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15;
dmux_1x16 dut(.i(i),.s0(s0),.s1(s1),.s2(s2),.s3(s3),.y0(y0),.y1(y1),.y2(y2),.y3(y3),.y4(y4),.y5(y5),.y6(y6),.y7(y7),.y8(y8),.y9(y9),.y10(y10),.y11(y11),.y12(y12),.y13(y13),.y14(y14),.y15(y15));
initial begin
	repeat(30)begin
	{i,s0,s1,s2,s3}=$random;
	#1;
$display("\t %0t i=%b || s3=%b  s2=%b  s1=%b  s0=%b || y0=%b  y1=%b  y2=%b  y3=%b  y4=%b  y5=%b  y6=%b  y7=%b  y8=%b  y9=%b  y10=%b  y11=%b  y12=%b  y13=%b  y14=%b  y15=%b",$time,i,s3,s2,s1,s0,y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15);
	end
	end
endmodule
*/

/*
output
 1 i=0  || s3=0  s2=0  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 2 i=0  || s3=1  s2=0  s1=0  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 3 i=0  || s3=1  s2=0  s1=0  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 4 i=0  || s3=1  s2=1  s1=0  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 5 i=0  || s3=1  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 6 i=0  || s3=1  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 7 i=0  || s3=1  s2=0  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 8 i=1  || s3=0  s2=1  s1=0  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=1  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 9 i=0  || s3=1  s2=0  s1=0  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 10 i=0 || s3=1  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 11 i=1 || s3=0  s2=1  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=1  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 12 i=1 || s3=1  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=1  y12=0  y13=0  y14=0  y15=0
 13 i=0 || s3=1  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 14 i=0 || s3=0  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 15 i=1 || s3=1  s2=0  s1=0  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=1  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 16 i=0 || s3=0  s2=1  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 17 i=0 || s3=1  s2=0  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 18 i=0 || s3=0  s2=1  s1=0  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 19 i=0 || s3=1  s2=0  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 20 i=1 || s3=1  s2=1  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=1  y15=0
 21 i=1 || s3=0  s2=1  s1=0  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=1  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 22 i=0 || s3=1  s2=1  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 23 i=1 || s3=0  s2=1  s1=0  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=1  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 24 i=0 || s3=0  s2=1  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 25 i=0 || s3=0  s2=0  s1=0  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 26 i=0 || s3=1  s2=0  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 27 i=1 || s3=0  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=1  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 28 i=1 || s3=1  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=1  y12=0  y13=0  y14=0  y15=0
 29 i=0 || s3=1  s2=0  s1=1  s0=1 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
 30 i=0 || s3=1  s2=0  s1=1  s0=0 || y0=0  y1=0  y2=0  y3=0  y4=0  y5=0  y6=0  y7=0  y8=0  y9=0  y10=0  y11=0  y12=0  y13=0  y14=0  y15=0
*/
